library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity LUT_32_16 is
    Port ( D : in STD_LOGIC_VECTOR (4 downto 0);
           I : out STD_LOGIC_VECTOR (15 downto 0));
end LUT_32_16;

architecture Behavioral of LUT_32_16 is
    type rom_type is array (0 to 31) of std_logic_vector(15 downto 0);
        signal Instruction_ROM : rom_type :=(
           "0010111000000001",
           "0010001000000101",
           "0010010000000001",
           "0001010000000000",
           "0101111001000000",
           "0000001010000000",
           "0011001000000110",
           "0011000000000100",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000", 
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000",
           "0000000000000000"  
        );  
begin
    I <= Instruction_ROM(to_integer(unsigned(D)));
end Behavioral;
