library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Nanoprocessor is
end Nanoprocessor;

architecture Behavioral of Nanoprocessor is

begin


end Behavioral;
