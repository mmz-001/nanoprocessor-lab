library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Frame_LUT is
    Port ( D : in STD_LOGIC_VECTOR (7 downto 0);
           Seg_Out_0 : out STD_LOGIC_VECTOR (7 downto 0);
           Seg_Out_1 : out STD_LOGIC_VECTOR (7 downto 0);
           Seg_Out_2 : out STD_LOGIC_VECTOR (7 downto 0);
           Seg_Out_3 : out STD_LOGIC_VECTOR (7 downto 0));
end Frame_LUT;

architecture Behavioral of Frame_LUT is
    signal I : STD_LOGIC_VECTOR (31 downto 0);
    signal I_Wire : STD_LOGIC_VECTOR (31 downto 0);
    
    type rom_type is array (0 to 255) of std_logic_vector(31 downto 0);
        signal Frame_ROM : rom_type :=(
            "11111111111111111111111111111111",
            "11011111111111111111111111111111",
            "11001111111111111111111111111111",
            "11000111111111111111111111111111",
            "01100111111101111111111111111111",
            "01110111011101111111011111111111",
            "11111111011101110111011111110111",
            "11111111111111110111011111110011",
            "11111111111111111111111111110001",
            "11111111111111111111111111111000",
            "11111111111111111111111011111100",
            "11111111111111101111111011111110",
            "11111110111111101111111011111111",
            "11011110111111101111111111111111",
            "11001110111111111111111111111111",
            "11000111111111111111111111111111",
            "01100111111101111111111111111111",
            "01110111011101111111011111111111",
            "11111111011101110111011111110111",
            "11111111111111110111011111110011",
            "11111111111111111111111111110001",
            "11111111111111111111111111111000",
            "11111111111111111111111011111100",
            "11111111111111101111111011111110",
            "11111110111111101111111011111111",
            "11011110111111101111111111111111",
            "11001110111111111111111111111111",
            "11000111111111111111111111111111",
            "01100111111101111111111111111111",
            "01110111011101111111011111111111",
            "11111111011101110111011111110111",
            "11111111111111110111011111110011",
            "11111111111111111111111111110001",
            "11111111111111111111111111111000",
            "11111111111111111111111011111100",
            "11111111111111101111111011111110",
            "11111110111111101111111011111111",
            "11011110111111101111111111111111",
            "11001110111111111111111111111111",
            "11000111111111111111111111111111",
            "01100111111101111111111111111111",
            "01110111011101111111011111111111",
            "11111111011101110111011111110111",
            "11111111111111110111011111110011",
            "11111111111111111111111111110001",
            "11111111111111111111111111111000",
            "11111111111111111111111011111100",
            "11111111111111101111111011111110",
            "11111110111111101111111011111111",
            "11011110111111101111111111111111",
            "11001110111111111111111111111111",
            "11001111111111111111111111111111",
            "11101111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "10001000111111111111111111111111",
            "10000011111111111111111111111111",
            "10100001111111111111111111111111",
            "10110000111111111111111111111111",
            "11110001111111111111111111111111",
            "10001100111111111111111111111111",
            "10011000111111111111111111111111",
            "11011000111111111111111111111111",
            "11100011111111111111111111111111",
            "10010010111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110111111111111111111111111",
            "11000110100010011111111111111111",
            "11000110100001101111111111111111",
            "11000110110001111111111111111111",
            "11000110110001111111111111111111",
            "11000110110000001111111111111111",
            "11000110100011101111111111111111",
            "11000110110011101111111111111111",
            "11000110110011111111111111111111",
            "11000110100001101111111111111111",
            "11000110101010111111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101111111111111111",
            "11000110100100101010000111111111",
            "11000110100100101111100111111111",
            "11000110100100101100001011111111",
            "11000110100100101111100111111111",
            "11000110100100101000011111111111",
            "11000110100100101000100011111111",
            "11000110100100101100011111111111",
            "11000110100100101111100111111111",
            "11000110100100101010010011111111",
            "11000110100100101011000011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000110100100101000011011111111",
            "11000111100100101000011011111111",
            "11100111100100101000011011111111",
            "11110111100100101000011011111111",
            "11111111100100101000011011111111",
            "11111111100100111000011011111111",
            "11111111101100111000011011111111",
            "11111111111100111000011011111111",
            "11111111111101111000011011111111",
            "11111111111111111000011011111111",
            "11111111111111111000011111111111",
            "11111111111111111010011111111111",
            "11111111111111111110011111111111",
            "11111111111111111111011111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111101111111111111111",
            "11111111100111011111111111111111",
            "11111111110000001111111111111111",
            "11111111110000001111111111111111",
            "11111111110000001111111111111111",
            "11111111110000001111111111111111",
            "11111110110000001111111111111111",
            "10011110110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "10100100110000001111111111111111",
            "11111111101001001100000011111111",
            "11111111111111111010010011000000",
            "11111111111111111111111110100100",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111",
            "11111111111111111111111111111111"            
        );  
begin
    I_Wire <= Frame_ROM(to_integer(unsigned(D)));
    I <= I_Wire;
    Seg_Out_0 <= I_Wire(7 downto 0);
    Seg_Out_1 <= I_Wire(15 downto 8);
    Seg_Out_2 <= I_Wire(23 downto 16);
    Seg_Out_3 <= I_Wire(31 downto 24);
end Behavioral;
