library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Ins_Decoder_16_TB is

end Ins_Decoder_16_TB;

architecture Behavioral of Ins_Decoder_16_TB is
component Ins_Decoder_16
  Port (
    I : in STD_LOGIC_VECTOR (15 downto 0); -- 16 bit instruction
    R_In : in STD_LOGIC_VECTOR (7 downto 0);  -- Input Register
    Zero, Overflow, Negative, Interrupt : in STD_LOGIC;
    R_En, RA_Sel, RB_Sel : out STD_LOGIC_VECTOR (2 downto 0);
    Jmp_Flag : out STD_LOGIC;
    AU_Sel: out STD_LOGIC_VECTOR (2 downto 0);
    Load_Sel : out STD_LOGIC_VECTOR ( 1 downto 0);
    Jmp_Addr : out STD_LOGIC_VECTOR (4 downto 0);
    Im_Val : out STD_LOGIC_VECTOR (7 downto 0));
end component;

Signal I : STD_LOGIC_VECTOR (15 downto 0); -- 16 bit instruction
Signal R_In : STD_LOGIC_VECTOR (7 downto 0);  -- Input Register
Signal Zero, Overflow, Negative, Interrupt : STD_LOGIC;
Signal R_En, RA_Sel, RB_Sel : STD_LOGIC_VECTOR (2 downto 0);
Signal Jmp_Flag : STD_LOGIC;
Signal AU_Sel: STD_LOGIC_VECTOR (2 downto 0);
Signal Load_Sel : STD_LOGIC_VECTOR ( 1 downto 0);
Signal Jmp_Addr : STD_LOGIC_VECTOR (4 downto 0);
Signal Im_Val : STD_LOGIC_VECTOR (7 downto 0);

begin
UUT: Ins_Decoder_16
port map(
    I => I,
    R_In =>R_In,
    Zero =>Zero,
    Overflow =>Overflow,
    Negative =>Negative,
    Interrupt =>Interrupt,
    R_En => R_En,
    RA_Sel => RA_Sel,
    RB_Sel => RB_Sel,
    JMP_Flag => Jmp_Flag,
    AU_Sel => AU_Sel,
    Load_Sel => Load_Sel,
    Jmp_Addr => Jmp_Addr,
    Im_Val => Im_Val);

process
begin
-- MOVI, register 8 (111), value = 10 (00001010)
I <= "0010111000001010";
wait for 100 ns;
end process;

end Behavioral;
